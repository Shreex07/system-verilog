`timescale 1ns / 1ps


module NOTgate(input logic a,
    output logic y
    );
assign y = ~a;
endmodule
